/*
  Jonathan Joslin 7/12/25
  WriteToCache module writes data from CPU registers to a selected cache way in a set-associative cache.
  - NUM_WAYS: Number of cache ways (default 4).
  - DATA_WIDTH: Width of data bus (default 32 bits).
  - OFFSET_WIDTH: Width of offset field for addressing within a cache line.
  - Interfaces: Connects to WayInterface (cache ways) and WriteToCacheInterface (CPU write requests).
  - Assumes synchronous operation with active-low reset.
  - Decoupled from control module
*/
module WriteToCache #(
  parameter int NUM_WAYS    = 4,
  parameter int DATA_WIDTH  = 32,
  parameter int OFFSET_WIDTH
)(
  input logic                 clk, reset_n,
  WayInterface.write          wayIfs[NUM_WAYS],
  WriteToCacheInterface.slave writeToCacheIf
);

  // Data registers to latch the write request, decoupling from the control module.
  logic [NUM_WAYS - 1:0]      target_one_hot;
  logic [OFFSET_WIDTH - 1:0]  w_offset;
  logic [DATA_WIDTH - 1:0]    w_data; 
  logic [2:0]                 w_id;             // ID used by the controller to detemine if write request was started 
  
  // ----------------------------------------
  // Sending
  // ----------------------------------------
  // One-hot encoding to send data to correct way
  generate
    for(genvar i = 0; i < NUM_WAYS; i++) begin
      assign wayIfs[i].offset = w_offset;
      assign wayIfs[i].w_en   = (w_state == WAIT_FOR_ACK) & target_one_hot[i];
      assign wayIfs[i].dataIn = w_data;
    end
  endgenerate

  // ----------------------------------------
  // Receiving 
  // ----------------------------------------
  logic                   w_ack;
  logic [NUM_WAYS - 1:0]  ack_buffer;

  // Collect write acknowledgments from all ways
  generate
    for(genvar i = 0; i < NUM_WAYS; i++) begin
      assign ack_buffer[i] = wayIfs[i].w_ack;
    end
  endgenerate


  // A single acknowledgement signal is generated by OR-ing all individual acks.
  // This assumes only the way that was written to will assert its w_ack.
  assign w_ack = |ack_buffer;
  

  // ----------------------------------------
  // Flow Control 
  // ----------------------------------------
 
  typedef enum logic [0:0] { 
    IDLE,
    WAIT_FOR_ACK
  } w_state_t;

  w_state_t w_state;

  // Ready to recieve new request when in IDLE
  assign writeToCacheIf.ready         = w_state == IDLE;  

  // The ID of the transaction currently being processed.
  assign writeToCacheIf.id_in_progress = w_id;

  // This process manages the write transaction, latching data and generating control signals.
  always_ff @(posedge clk or negedge reset_n) begin
    if(!reset_n) begin
      w_state             <= IDLE;
      target_one_hot      <= '0;
      w_offset            <= '0;
      w_data              <= '0;
      w_id                <= '0;
    end
    else begin
      case(w_state)
        IDLE : begin
          if(writeToCacheIf.request) begin
            w_state         <= WAIT_FOR_ACK;
            w_offset        <= writeToCacheIf.offset;
            w_data          <= writeToCacheIf.w_data;
            target_one_hot  <= writeToCacheIf.targetWay;
            w_id            <= writeToCacheIf.write_id;
          end
        end
        WAIT_FOR_ACK : begin
          if(w_ack) begin
            w_state             <= IDLE;
            target_one_hot      <= '0;
            w_offset            <= '0;
            w_data              <= '0;
          end
        end
        default: begin
          w_state             <= IDLE;
          target_one_hot      <= '0;
          w_offset            <= '0;
          w_data              <= '0;
        end
      endcase
    end
  end






endmodule